`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:47:24 12/10/2016 
// Design Name: 
// Module Name:    Sixty_Four_Bit_Sign_Extender 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Sixty_Four_Bit_Sign_Extender(
	input signed [6:0] in,
	output signed [63:0] out
    ); 
 assign out =in;

endmodule
